library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity tb_output_mux is
--  Port ( );
end tb_output_mux;

architecture Behavioral of tb_output_mux is

begin


end Behavioral;
